module background ( input [7:0]	addr,
						output [255:0]	data
					 );

	parameter ADDR_WIDTH = 8;
   parameter DATA_WIDTH =  256;
	logic [ADDR_WIDTH-1:0] addr_reg;

	// ROM definition
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {

256'b 0000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000,
256'b 0000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110,
256'b 0001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
256'b 0001000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001,
256'b 0011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000001111111111111111111111100000000000000000000000111111111111111111111111111111110000000000000000000010000000100000000000000000000011111111111111111111111111111111000000000000000000000011111111111111111111111000000000000000000001100,
256'b 0011001000000000000000000010000000000000000000000010000000000000000000001000000000000000000000000000000001000000000000000000010000000100000000000000000001100000000000000000000000000000000100000000000000000000100000000000000000000000100000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000010000000000000000000000000000000000100000000000000000011000000100000000000000000001000000000000000000000000000000000110000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000011000000000000000000000010000000000000000000001000000000000000000000000000000011000000000000000000001100011000000000000000000000100000000000000000000000000000001100000000000000000000110000000000000000000000100000000000000000001100,
256'b 0011001000000000000000000000111111111111111111111100000000000000000000000111111111111111111111111111111100000000000000000000000011110000000000000000000000011111111111111111111111111111110000000000000000000000001111111111111111111111000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000001111111111111111111111100000000000000000000000111100000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000000011111000000000000000000000011111111111111111111111000000000000000000001100,
256'b 0011001000000000000000000010000000000000000000000010000000000000000000001000011000000000000000000001000000000000000000000000000000000000000000000000000000000001100000000000000000000100000100000000000000000000100000000000000000000000100000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000010000000000000000000000011000000000000000000110000001100000000000000000001000000000000000000000000000000000000000000000000000000000001100000000000000000001000000010000000000000000000100000000000000000000000110000000000000000001100,
256'b 0011001000000000000000000001111111111111111111111100000000000000000000110000001100000000000000000000111111111111111111111111000000000000111111111111111111111111000000000000000000001000000010000000000000000000011111111111111111111111000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000100000000011000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000000100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011000100000000000000000000000000000000000000000000000000000000000000110000000010000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000110000000010000000000000000000000000000000000000000000000000000000000000010000,
256'b 0001100011111111111111111111111111111111111111111110000000000000000000110000000001111111111111111111111110000000000000000000010000000100000000000000000000111111111111111111111111000000000010000000000000000000011111111111111111111111111111111111111111100001,
256'b 0000111000000000000000000000000000000000000000000001000000000000000000110000000000000000000000000000000001100000000000000000010000000100000000000000000001000000000000000000000000000000000010000000000000000001100000000000000000000000000000000000000000000111,
256'b 0000001111111111111111111111111111111111111111110001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000011111111111111111111111111111111111111111000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000000000000000000000000000000001000000000000000000001000001000000000000000000000100000000000000000000000000000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000000001111111111111111111111110000000000000000000000111110000000000000000000000011111111111111111111111100000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000011111111111111111111110000000000000000000111111111111111111111100000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000010000000000000000000011111111111111111111100000000000000000000110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000010000000000000000000011111111111111111111100000000000000000000110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000010011111111111111111111000000000000000001111111111111111111100110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0011111111111111111111111111111111111111111111110001000000000000000000110000001100000000000000000010011000000000000000000000000000000000000000000000000000000100110000000000000000001000000010000000000000000001000011111111111111111111111111111111111111111111,
256'b 0000000000000000000000000000000000000000000000000001000000000000000000010000001100000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000001000000010000000000000000001000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000010000000000000000000001000010000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000100001100000000000000000000110000000000000000000000000000000000000000000000,
256'b 0001111111111111111111111111111111111111111111111100000000000000000000000111100000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000011110000000000000000000000001111111111111111111111111111111111111111111111,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
256'b 0011111111111111111111111111111111111111111111111100000000000000000000000111100000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000011111000000000000000000000011111111111111111111111111111111111111111111111,
256'b 0000000000000000000000000000000000000000000000000010000000000000000000001000011000000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000000100000100000000000000000000100000000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000000001000000000000000000110000001100000000000000000010010000000000000000000000000000000000000000000000000000000100110000000000000000001000000010000000000000000001000000000000000000000000000000000000000000000000,
256'b 0011111111111111111111111111111111111111111111110001000000000000000000110000001100000000000000000010011000000000000000000000000000000000000000000000000000001100110000000000000000001000000010000000000000000001000111111111111111111111111111111111111111111111,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000010001111111111111111111111111111111111111111111111111111111100110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000011000000000000000000000000000000000000000000000000000000000000100000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000000000000000000000000000000000000000000001001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001001100000000000000000000000000000000000000000000,
256'b 0000000111111111111111111111111111111111111111110001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000111111111111111111111111111111111111111110000,
256'b 0000011000000000000000000000000000000000000000000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000000000000000000000000000000000000000001110,
256'b 0001100000000000000000000000000000000000000000000010000000000000000000001000011000000000000000000001000000000000000000000000000000000000000000000000000000000001100000000000000000000100000100000000000000000000100000000000000000000000000000000000000000000001,
256'b 0001100011111111111111111111111111111111111111111100000000000000000000000111100000000000000000000000111111111111111111111111000000000001111111111111111111111110000000000000000000000011111000000000000000000000011111111111111111111111111111111111111111110001,
256'b 0011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000001111111111111111111111100000000000000000000000111111111111111111111111111111100000000000000000000010000000100000000000000000000011111111111111111111111111111110000000000000000000000001111111111111111111111000000000000000000001100,
256'b 0011001000000000000000000011000000000000000000000010000000000000000000001000000000000000000000000000000011000000000000000000010000000100000000000000000000100000000000000000000000000000001100000000000000000000110000000000000000000000100000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000010000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000110000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000001000000000000000000010000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000010000000000000000001000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000011000000000000000000000001000000000000000000001000000000000000000000000000000011000000000000000000001100001000000000000000000000100000000000000000000000000000001100000000000000000001000000000000000000000000100000000000000000001100,
256'b 0011001000000000000000000000111111111111111000000001000000000000000000000111111111111111111111111111111100000000000000000000000011110000000000000000000000011111111111111111111111111111110000000000000000000001000000000111111111111111000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000001100,
256'b 0011000100000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000011000,
256'b 0011000011111111111111100000000000000000000100000001000000000000000000000111100000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000000011111000000000000000000001000000010000000000000000000001111111111111100000,
256'b 0011000000000000000000010000000000000000000100000001000000000000000000001000011000000000000000000001000000000000000000000000000000000000000000000000000000000001100000000000000000000100000100000000000000000001000000010000000000000000000110000000000000000000,
256'b 0011000000000000000000001000000000000000000100000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000010000000000000000001100000000000000000000,
256'b 0011000000000000000000001000000000000000000100000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000010000000000000000001100000000000000000000,
256'b 0011000000000000000000001000000000000000000100000001000000000000000000110000001100000000000000000010000000000000000000000000000000000000000000000000000000000000110000000000000000001000000010000000000000000001000000010000000000000000001100000000000000000000,
256'b 0011000000000000000000010000000000000000000010000011000000000000000000110000001100000000000000000011000000000000000000000000000000000000000000000000000000000000100000000000000000001000000010000000000000000000100000110000000000000000000100000000000000000000,
256'b 0011000011111111111111100000000000000000000001111100000000000000000000110000001100000000000000000000111111111111111111111111000000000000111111111111111111111111000000000000000000001000000010000000000000000000011111000000000000000000000011111111111111100000,
256'b 0011000100000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000100000000011000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000011000,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000110000000100000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000110000000001000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000001111111111111111111111111111111111111111110000000000001111111111111111111111110000000000000000000010000000100000000000000000000111111111111111111111111000000000000111111111111111111111111111111111111111111100000000000000000001100,
256'b 0011001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000100000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001100,
256'b 0011001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001000001000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001100,
256'b 0011001000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
256'b 0011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000,
256'b 0001000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001,
256'b 0001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
256'b 0000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110,
256'b 0000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000
};

	assign data = ROM[addr];

endmodule 