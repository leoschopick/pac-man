module ghostfont ( input logic [4:0]	addr,
						output logic [31:0]	data
					 );

	parameter ADDR_WIDTH = 5;
   parameter DATA_WIDTH =  32;
	logic [ADDR_WIDTH-1:0] addr_reg;

	// ROM definition
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {

		//Pacman facing right
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000111111111110000000000,
		32'b 00000000011111111111111000000000,
		32'b 00000000111111111111111100000000,
		32'b 00000001111111111111111110000000,
		32'b 00000011111111111111111111000000,
		32'b 00000111111111111111111111100000,
		32'b 00000111110011111111100111100000,
		32'b 00001111100001111111000011110000,
		32'b 00001111100001111111000011110000,
		32'b 00001111100001111111000011110000,
		32'b 00011111110011111111100111111000,
		32'b 00011111111111111111111111111000,
		32'b 00011111111111111111111111111000,
		32'b 00011111111111111111111111111000,
		32'b 00011111111111111111111111111000,
		32'b 00011111111111111111111111111000,
		32'b 00011110111111110111111110111000,
		32'b 00011100011111100011111100011000,
		32'b 00011100001111100001111000011000,
		32'b 00011000000111000000111000011000,
		32'b 00010000000010000000010000001000,
		32'b 00010000000010000000010000001000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000,
		32'b 00000000000000000000000000000000

	};

	assign data = ROM[addr];

endmodule